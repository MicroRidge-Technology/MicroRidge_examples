`default_nettype none
/**/
`timescale 1ns/1ns
module dc_fifo
#(parameter type T)
(
 input logic clka;
 input logic clkb;
 input
);
endmodule
`default_nettype wire
